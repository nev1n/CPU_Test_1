
library ieee;
use ieee.std_logic_1164.all;

entity ADDER_TB is 
end ADDER_TB;

architecture behaviour_ADDER_TB of ADDER_TB is